--pacote de parametros do projeto
library ieee;
use ieee.std_logic_1164.all;

package parametros is

	--comprimento da janela de media movel
	constant Mbits : natural := 4;

	--comprimento da palavra
	constant Nbits : natural := 8;

end package parametros;

package body parametros is

end;
