library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package parametros is

	constant Kbits : natural := 4;

end package parametros;

package body parametros is

end;
